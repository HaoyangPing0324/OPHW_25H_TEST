//****************************************Copyright (c)***********************************//
//ԭ�Ӹ����߽�ѧƽ̨��www.yuanzige.com
//����֧�֣�www.openedv.com
//�Ա����̣�http://openedv.taobao.com 
//��ע΢�Ź���ƽ̨΢�źţ�"����ԭ��"����ѻ�ȡZYNQ & FPGA & STM32 & LINUX���ϡ�
//��Ȩ���У�����ؾ���
//Copyright(C) ����ԭ�� 2018-2028
//All rights reserved                                  
//----------------------------------------------------------------------------------------
// File name:           rgmii_tx
// Last modified Date:  2020/2/13 9:20:14
// Last Version:        V1.0
// Descriptions:        RGMII����ģ��
//----------------------------------------------------------------------------------------
// Created by:          ����ԭ��
// Created date:        2020/2/13 9:20:14
// Version:             V1.0
// Descriptions:        The original version
//
//----------------------------------------------------------------------------------------
//****************************************************************************************//

module rgmii_tx(
    //GMII���Ͷ˿�
    input              gmii_tx_clk , //GMII����ʱ��    
    input              gmii_tx_en  , //GMII���������Ч�ź�
    input       [7:0]  gmii_txd    , //GMII�������        
    
    //RGMII���Ͷ˿�
    output             rgmii_txc   , //RGMII��������ʱ��    
    output             rgmii_tx_ctl, //RGMII���������Ч�ź�
    output      [3:0]  rgmii_txd     //RGMII�������     
    );

//*****************************************************
//**                    main code
//*****************************************************

assign rgmii_txc = gmii_tx_clk;

//���˫�ز����Ĵ��� (rgmii_tx_ctl)

GTP_ODDR_E1 #(
    .GRS_EN("TRUE"),
    .ODDR_MODE("SAME_EDGE"),
    .RS_TYPE("SYNC_RESET") 
) u_ODDR_inst_tx_ctl (
    .Q(rgmii_tx_ctl),  // OUTPUT  
    .CE(1'b1), // INPUT  
    .CLK(gmii_tx_clk),// INPUT  
    .D0(gmii_tx_en), // INPUT  
    .D1(gmii_tx_en), // INPUT  
    .RS(1'b0)  // INPUT  
);

genvar i;
generate for (i=0; i<4; i=i+1)
    begin : txdata_bus
        //���˫�ز����Ĵ��� (rgmii_txd)

GTP_ODDR_E1 #(
    .GRS_EN("TRUE"),
    .ODDR_MODE("SAME_EDGE"),
    .RS_TYPE("SYNC_RESET") 
) u_ODDR_inst_txdata (
    .Q(rgmii_txd[i]),  // OUTPUT  
    .CE(1'b1), // INPUT  
    .CLK(gmii_tx_clk),// INPUT  
    .D0(gmii_txd[i]), // INPUT  
    .D1(gmii_txd[4+i]), // INPUT  
    .RS(1'b0)  // INPUT  
);       
    end
endgenerate

endmodule