//****************************************Copyright (c)***********************************//
//ԭ�Ӹ����߽�ѧƽ̨��www.yuanzige.com
//����֧�֣�www.openedv.com
//�Ա����̣�http://openedv.taobao.com 
//��ע΢�Ź���ƽ̨΢�źţ�"����ԭ��"����ѻ�ȡZYNQ & FPGA & STM32 & LINUX���ϡ�
//��Ȩ���У�����ؾ���
//Copyright(C) ����ԭ�� 2018-2028
//All rights reserved                                  
//----------------------------------------------------------------------------------------
// File name:           rgmii_rx
// Last modified Date:  2020/2/13 9:20:14
// Last Version:        V1.0
// Descriptions:        RGMII����ģ��
//----------------------------------------------------------------------------------------
// Created by:          ����ԭ��
// Created date:        2020/2/13 9:20:14
// Version:             V1.0
// Descriptions:        The original version
//
//----------------------------------------------------------------------------------------
//****************************************************************************************//

module rgmii_rx(
    input              idelay_clk  , //200Mhzʱ�ӣ�IDELAYʱ��
    
    //��̫��RGMII�ӿ�
    input              rgmii_rxc   , //RGMII����ʱ��
    input              rgmii_rx_ctl, //RGMII�������ݿ����ź�
    input       [3:0]  rgmii_rxd   , //RGMII��������    

    //��̫��GMII�ӿ�
    output             gmii_rx_clk , //GMII����ʱ��
    output             gmii_rx_dv  , //GMII����������Ч�ź�
    output      [7:0]  gmii_rxd      //GMII��������   
    );

//wire define
wire         rgmii_rxc_bufg;     //ȫ��ʱ�ӻ���
wire         rgmii_rxc_bufio;    //ȫ��ʱ��IO����
wire  [3:0]  rgmii_rxd_delay;    //rgmii_rxd������ʱ
wire         rgmii_rx_ctl_delay; //rgmii_rx_ctl������ʱ
wire  [1:0]  gmii_rxdv_t;        //��λGMII������Ч�ź� 

//*****************************************************
//**                    main code
//*****************************************************

assign gmii_rx_clk = rgmii_rxc_bufg;
assign gmii_rx_dv = gmii_rxdv_t[0] & gmii_rxdv_t[1];

//ȫ��ʱ�ӻ���
GTP_CLKBUFG BUFG_inst(
    .CLKOUT(rgmii_rxc_bufg),// OUTPUT  
    .CLKIN(rgmii_rxc)  // INPUT  
);

//ȫ��ʱ��IO����

GTP_IOCLKBUF #(
    .GATE_EN("FALSE") 
) u_GTP_IOCLKBUF (
    .CLKOUT(rgmii_rxc_bufio),// OUTPUT  
    .CLKIN(rgmii_rxc), // INPUT  
    .DI(1'b1)     // INPUT  
);

////����˫�ز����Ĵ���
GTP_IDDR_E1 #(
    .GRS_EN("TRUE"),
    .IDDR_MODE("SAME_PIPELINED"),
    .RS_TYPE(" SYNC_RESET") 
) u_iddr_rx_ctl (
    .Q0(gmii_rxdv_t[0]), // OUTPUT  
    .Q1(gmii_rxdv_t[1]), // OUTPUT  
    .CE(1'b1), // INPUT  
    .CLK(rgmii_rxc_bufio),// INPUT  
    .D(rgmii_rx_ctl),  // INPUT  
    .RS(1'b0)  // INPUT  
);

//rgmii_rxd������ʱ��˫�ز���
genvar i;
generate for (i=0; i<4; i=i+1) 
    begin : rxdata_bus	
GTP_IDDR_E1 #(
    .GRS_EN("TRUE"),
    .IDDR_MODE("SAME_PIPELINED"),
    .RS_TYPE(" SYNC_RESET") 
) u_iddr_rxd (
    .Q0(gmii_rxd[i]), // OUTPUT  
    .Q1(gmii_rxd[4+i]), // OUTPUT  
    .CE(1'b1), // INPUT  
    .CLK(rgmii_rxc_bufio),// INPUT  
    .D(rgmii_rxd[i]),  // INPUT  
    .RS(1'b0)  // INPUT  
);		
		
    end
endgenerate

endmodule