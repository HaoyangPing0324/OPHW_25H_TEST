`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//Copyright(C) ����ԭ�� 2023-2033
// Revised By HaoyangPing_PKU
//
//////////////////////////////////////////////////////////////////////////////////
`define UD #1
module video_display # (
    parameter                            COCLOR_DEPP=8, // number of bits per channel
    parameter                            X_BITS=12,
    parameter                            Y_BITS=12,
    parameter                            H_ACT = 12'd1280,
    parameter                            V_ACT = 12'd720
)(                                       
    input                                rstn, 
    input                                pix_clk,
    input [X_BITS-1:0]                   act_x,
	input [Y_BITS-1:0]                   act_y,
    input                                vs_in, 
    input                                hs_in, 
    input                                de_in,
    
    output reg                           vs_out, 
    output reg                           hs_out, 
    output reg                           de_out,
    output reg [3*COCLOR_DEPP-1:0]       pixel_data 
);
    
    always @(posedge pix_clk)
    begin
        vs_out <= `UD vs_in;
        hs_out <= `UD hs_in;
        de_out <= `UD de_in;
    end

//parameter define    
parameter  DIV_CNT = 22'd750000;				//��Ƶ������

localparam SIDE_W  = 11'd40;                    //��Ļ�߿���
localparam BLOCK_W = 11'd40;                    //������
localparam BLUE    = 24'h0000ff;    			//��Ļ�߿���ɫ ��ɫ
localparam WHITE   = 24'hffffff;    			//������ɫ ��ɫ
localparam BLACK   = 24'h000000;    			//������ɫ ��ɫ


//reg define
reg [10:0] block_x = SIDE_W ;                   //�������ϽǺ�����
reg [10:0] block_y = SIDE_W ;                   //�������Ͻ�������
reg [21:0] div_cnt;                             //ʱ�ӷ�Ƶ������
reg        h_direct;                            //����ˮƽ�ƶ�����1�����ƣ�0������
reg        v_direct;                            //������ֱ�ƶ�����1�����£�0������

//wire define   
wire move_en;                                   //�����ƶ�ʹ���źţ�Ƶ��Ϊ100hz

//*****************************************************
//**                    main code
//*****************************************************
assign move_en = (div_cnt == DIV_CNT) ? 1'b1 : 1'b0;

//ͨ����div����ʱ�Ӽ�����ʵ��ʱ�ӷ�Ƶ
always @(posedge pix_clk or negedge rstn) begin         
    if (!rstn)
        div_cnt <= 22'd0;
    else begin
        if(div_cnt < DIV_CNT) 
            div_cnt <= div_cnt + 1'b1;
        else
            div_cnt <= 22'd0;                   //������10ms������
    end
end

//�������ƶ����߽�ʱ���ı��ƶ�����
always @(posedge pix_clk or negedge rstn) begin         
    if (!rstn) begin
        h_direct <= 1'b1;                       //�����ʼˮƽ�����ƶ�
        v_direct <= 1'b1;                       //�����ʼ��ֱ�����ƶ�
    end
    else begin
        if(block_x == SIDE_W + 1'b1)            //������߽�ʱ��ˮƽ����
            h_direct <= 1'b1;               
        else                                    //�����ұ߽�ʱ��ˮƽ����
        if(block_x == H_ACT - SIDE_W - BLOCK_W + 1'b1)
            h_direct <= 1'b0;               
        else
            h_direct <= h_direct;
            
        if(block_y == SIDE_W + 1'b1)            //�����ϱ߽�ʱ����ֱ����
            v_direct <= 1'b1;                
        else                                    //�����±߽�ʱ����ֱ����
        if(block_y == V_ACT - SIDE_W - BLOCK_W + 1'b1)
            v_direct <= 1'b0;               
        else
            v_direct <= v_direct;
    end
end

//���ݷ����ƶ����򣬸ı����ݺ�����
always @(posedge pix_clk or negedge rstn) begin         
    if (!rstn) begin
        block_x <= SIDE_W + 1'b1;                     //�����ʼλ�ú�����
        block_y <= SIDE_W + 1'b1;                     //�����ʼλ��������
    end
    else if(move_en) begin
        if(h_direct) 
            block_x <= block_x + 1'b1;          //���������ƶ�
        else
            block_x <= block_x - 1'b1;          //���������ƶ�
            
        if(v_direct) 
            block_y <= block_y + 1'b1;          //���������ƶ�
        else
            block_y <= block_y - 1'b1;          //���������ƶ�
    end
    else begin
        block_x <= block_x;
        block_y <= block_y;
    end
end

//����ͬ��������Ʋ�ͬ����ɫ
always @(posedge pix_clk or negedge rstn) begin         
    if (!rstn) 
        pixel_data <= BLACK;
    else begin
        if(  (act_x < SIDE_W) || (act_x >= H_ACT - SIDE_W)
          || (act_y <= SIDE_W) || (act_y > V_ACT - SIDE_W))
            pixel_data <= BLUE;                 //������Ļ�߿�Ϊ��ɫ
        else
        if(  (act_x >= block_x - 1'b1) && (act_x < block_x + BLOCK_W - 1'b1)
          && (act_y >= block_y) && (act_y < block_y + BLOCK_W))
            pixel_data <= BLACK;                //���Ʒ���Ϊ��ɫ
        else
            pixel_data <= WHITE;                //���Ʊ���Ϊ��ɫ
    end
end

endmodule 