//gamma_table
module gamma_lookuptable
(
   input		[7:0]	video_data,
   output		reg[7:0]	gamma_data
);

always@(*)
begin
	case(video_data)
	8'd0 : gamma_data = 8'd0; 
	8'd1 : gamma_data = 8'd128; 
	8'd2 : gamma_data = 8'd139; 
	8'd3 : gamma_data = 8'd146; 
	8'd4 : gamma_data = 8'd152; 
	8'd5 : gamma_data = 8'd156; 
	8'd6 : gamma_data = 8'd160; 
	8'd7 : gamma_data = 8'd163; 
	8'd8 : gamma_data = 8'd165; 
	8'd9 : gamma_data = 8'd168; 
	8'd10 : gamma_data = 8'd170; 
	8'd11 : gamma_data = 8'd172; 
	8'd12 : gamma_data = 8'd174; 
	8'd13 : gamma_data = 8'd176; 
	8'd14 : gamma_data = 8'd177; 
	8'd15 : gamma_data = 8'd179; 
	8'd16 : gamma_data = 8'd180; 
	8'd17 : gamma_data = 8'd182; 
	8'd18 : gamma_data = 8'd183; 
	8'd19 : gamma_data = 8'd184; 
	8'd20 : gamma_data = 8'd186; 
	8'd21 : gamma_data = 8'd187; 
	8'd22 : gamma_data = 8'd188; 
	8'd23 : gamma_data = 8'd189; 
	8'd24 : gamma_data = 8'd190; 
	8'd25 : gamma_data = 8'd191; 
	8'd26 : gamma_data = 8'd192; 
	8'd27 : gamma_data = 8'd193; 
	8'd28 : gamma_data = 8'd193; 
	8'd29 : gamma_data = 8'd194; 
	8'd30 : gamma_data = 8'd195; 
	8'd31 : gamma_data = 8'd196; 
	8'd32 : gamma_data = 8'd197; 
	8'd33 : gamma_data = 8'd197; 
	8'd34 : gamma_data = 8'd198; 
	8'd35 : gamma_data = 8'd199; 
	8'd36 : gamma_data = 8'd200; 
	8'd37 : gamma_data = 8'd200; 
	8'd38 : gamma_data = 8'd201; 
	8'd39 : gamma_data = 8'd202; 
	8'd40 : gamma_data = 8'd202; 
	8'd41 : gamma_data = 8'd203; 
	8'd42 : gamma_data = 8'd204; 
	8'd43 : gamma_data = 8'd204; 
	8'd44 : gamma_data = 8'd205; 
	8'd45 : gamma_data = 8'd205; 
	8'd46 : gamma_data = 8'd206; 
	8'd47 : gamma_data = 8'd206; 
	8'd48 : gamma_data = 8'd207; 
	8'd49 : gamma_data = 8'd207; 
	8'd50 : gamma_data = 8'd208; 
	8'd51 : gamma_data = 8'd209; 
	8'd52 : gamma_data = 8'd209; 
	8'd53 : gamma_data = 8'd210; 
	8'd54 : gamma_data = 8'd210; 
	8'd55 : gamma_data = 8'd211; 
	8'd56 : gamma_data = 8'd211; 
	8'd57 : gamma_data = 8'd211; 
	8'd58 : gamma_data = 8'd212; 
	8'd59 : gamma_data = 8'd212; 
	8'd60 : gamma_data = 8'd213; 
	8'd61 : gamma_data = 8'd213; 
	8'd62 : gamma_data = 8'd214; 
	8'd63 : gamma_data = 8'd214; 
	8'd64 : gamma_data = 8'd215; 
	8'd65 : gamma_data = 8'd215; 
	8'd66 : gamma_data = 8'd215; 
	8'd67 : gamma_data = 8'd216; 
	8'd68 : gamma_data = 8'd216; 
	8'd69 : gamma_data = 8'd217; 
	8'd70 : gamma_data = 8'd217; 
	8'd71 : gamma_data = 8'd217; 
	8'd72 : gamma_data = 8'd218; 
	8'd73 : gamma_data = 8'd218; 
	8'd74 : gamma_data = 8'd218; 
	8'd75 : gamma_data = 8'd219; 
	8'd76 : gamma_data = 8'd219; 
	8'd77 : gamma_data = 8'd220; 
	8'd78 : gamma_data = 8'd220; 
	8'd79 : gamma_data = 8'd220; 
	8'd80 : gamma_data = 8'd221; 
	8'd81 : gamma_data = 8'd221; 
	8'd82 : gamma_data = 8'd221; 
	8'd83 : gamma_data = 8'd222; 
	8'd84 : gamma_data = 8'd222; 
	8'd85 : gamma_data = 8'd222; 
	8'd86 : gamma_data = 8'd223; 
	8'd87 : gamma_data = 8'd223; 
	8'd88 : gamma_data = 8'd223; 
	8'd89 : gamma_data = 8'd224; 
	8'd90 : gamma_data = 8'd224; 
	8'd91 : gamma_data = 8'd224; 
	8'd92 : gamma_data = 8'd224; 
	8'd93 : gamma_data = 8'd225; 
	8'd94 : gamma_data = 8'd225; 
	8'd95 : gamma_data = 8'd225; 
	8'd96 : gamma_data = 8'd226; 
	8'd97 : gamma_data = 8'd226; 
	8'd98 : gamma_data = 8'd226; 
	8'd99 : gamma_data = 8'd227; 
	8'd100 : gamma_data = 8'd227; 
	8'd101 : gamma_data = 8'd227; 
	8'd102 : gamma_data = 8'd227; 
	8'd103 : gamma_data = 8'd228; 
	8'd104 : gamma_data = 8'd228; 
	8'd105 : gamma_data = 8'd228; 
	8'd106 : gamma_data = 8'd228; 
	8'd107 : gamma_data = 8'd229; 
	8'd108 : gamma_data = 8'd229; 
	8'd109 : gamma_data = 8'd229; 
	8'd110 : gamma_data = 8'd230; 
	8'd111 : gamma_data = 8'd230; 
	8'd112 : gamma_data = 8'd230; 
	8'd113 : gamma_data = 8'd230; 
	8'd114 : gamma_data = 8'd231; 
	8'd115 : gamma_data = 8'd231; 
	8'd116 : gamma_data = 8'd231; 
	8'd117 : gamma_data = 8'd231; 
	8'd118 : gamma_data = 8'd232; 
	8'd119 : gamma_data = 8'd232; 
	8'd120 : gamma_data = 8'd232; 
	8'd121 : gamma_data = 8'd232; 
	8'd122 : gamma_data = 8'd233; 
	8'd123 : gamma_data = 8'd233; 
	8'd124 : gamma_data = 8'd233; 
	8'd125 : gamma_data = 8'd233; 
	8'd126 : gamma_data = 8'd233; 
	8'd127 : gamma_data = 8'd234; 
	8'd128 : gamma_data = 8'd234; 
	8'd129 : gamma_data = 8'd234; 
	8'd130 : gamma_data = 8'd234; 
	8'd131 : gamma_data = 8'd235; 
	8'd132 : gamma_data = 8'd235; 
	8'd133 : gamma_data = 8'd235; 
	8'd134 : gamma_data = 8'd235; 
	8'd135 : gamma_data = 8'd236; 
	8'd136 : gamma_data = 8'd236; 
	8'd137 : gamma_data = 8'd236; 
	8'd138 : gamma_data = 8'd236; 
	8'd139 : gamma_data = 8'd236; 
	8'd140 : gamma_data = 8'd237; 
	8'd141 : gamma_data = 8'd237; 
	8'd142 : gamma_data = 8'd237; 
	8'd143 : gamma_data = 8'd237; 
	8'd144 : gamma_data = 8'd237; 
	8'd145 : gamma_data = 8'd238; 
	8'd146 : gamma_data = 8'd238; 
	8'd147 : gamma_data = 8'd238; 
	8'd148 : gamma_data = 8'd238; 
	8'd149 : gamma_data = 8'd238; 
	8'd150 : gamma_data = 8'd239; 
	8'd151 : gamma_data = 8'd239; 
	8'd152 : gamma_data = 8'd239; 
	8'd153 : gamma_data = 8'd239; 
	8'd154 : gamma_data = 8'd239; 
	8'd155 : gamma_data = 8'd240; 
	8'd156 : gamma_data = 8'd240; 
	8'd157 : gamma_data = 8'd240; 
	8'd158 : gamma_data = 8'd240; 
	8'd159 : gamma_data = 8'd240; 
	8'd160 : gamma_data = 8'd241; 
	8'd161 : gamma_data = 8'd241; 
	8'd162 : gamma_data = 8'd241; 
	8'd163 : gamma_data = 8'd241; 
	8'd164 : gamma_data = 8'd241; 
	8'd165 : gamma_data = 8'd241; 
	8'd166 : gamma_data = 8'd242; 
	8'd167 : gamma_data = 8'd242; 
	8'd168 : gamma_data = 8'd242; 
	8'd169 : gamma_data = 8'd242; 
	8'd170 : gamma_data = 8'd242; 
	8'd171 : gamma_data = 8'd243; 
	8'd172 : gamma_data = 8'd243; 
	8'd173 : gamma_data = 8'd243; 
	8'd174 : gamma_data = 8'd243; 
	8'd175 : gamma_data = 8'd243; 
	8'd176 : gamma_data = 8'd243; 
	8'd177 : gamma_data = 8'd244; 
	8'd178 : gamma_data = 8'd244; 
	8'd179 : gamma_data = 8'd244; 
	8'd180 : gamma_data = 8'd244; 
	8'd181 : gamma_data = 8'd244; 
	8'd182 : gamma_data = 8'd244; 
	8'd183 : gamma_data = 8'd245; 
	8'd184 : gamma_data = 8'd245; 
	8'd185 : gamma_data = 8'd245; 
	8'd186 : gamma_data = 8'd245; 
	8'd187 : gamma_data = 8'd245; 
	8'd188 : gamma_data = 8'd245; 
	8'd189 : gamma_data = 8'd246; 
	8'd190 : gamma_data = 8'd246; 
	8'd191 : gamma_data = 8'd246; 
	8'd192 : gamma_data = 8'd246; 
	8'd193 : gamma_data = 8'd246; 
	8'd194 : gamma_data = 8'd246; 
	8'd195 : gamma_data = 8'd247; 
	8'd196 : gamma_data = 8'd247; 
	8'd197 : gamma_data = 8'd247; 
	8'd198 : gamma_data = 8'd247; 
	8'd199 : gamma_data = 8'd247; 
	8'd200 : gamma_data = 8'd247; 
	8'd201 : gamma_data = 8'd248; 
	8'd202 : gamma_data = 8'd248; 
	8'd203 : gamma_data = 8'd248; 
	8'd204 : gamma_data = 8'd248; 
	8'd205 : gamma_data = 8'd248; 
	8'd206 : gamma_data = 8'd248; 
	8'd207 : gamma_data = 8'd248; 
	8'd208 : gamma_data = 8'd249; 
	8'd209 : gamma_data = 8'd249; 
	8'd210 : gamma_data = 8'd249; 
	8'd211 : gamma_data = 8'd249; 
	8'd212 : gamma_data = 8'd249; 
	8'd213 : gamma_data = 8'd249; 
	8'd214 : gamma_data = 8'd249; 
	8'd215 : gamma_data = 8'd250; 
	8'd216 : gamma_data = 8'd250; 
	8'd217 : gamma_data = 8'd250; 
	8'd218 : gamma_data = 8'd250; 
	8'd219 : gamma_data = 8'd250; 
	8'd220 : gamma_data = 8'd250; 
	8'd221 : gamma_data = 8'd250; 
	8'd222 : gamma_data = 8'd251; 
	8'd223 : gamma_data = 8'd251; 
	8'd224 : gamma_data = 8'd251; 
	8'd225 : gamma_data = 8'd251; 
	8'd226 : gamma_data = 8'd251; 
	8'd227 : gamma_data = 8'd251; 
	8'd228 : gamma_data = 8'd251; 
	8'd229 : gamma_data = 8'd252; 
	8'd230 : gamma_data = 8'd252; 
	8'd231 : gamma_data = 8'd252; 
	8'd232 : gamma_data = 8'd252; 
	8'd233 : gamma_data = 8'd252; 
	8'd234 : gamma_data = 8'd252; 
	8'd235 : gamma_data = 8'd252; 
	8'd236 : gamma_data = 8'd253; 
	8'd237 : gamma_data = 8'd253; 
	8'd238 : gamma_data = 8'd253; 
	8'd239 : gamma_data = 8'd253; 
	8'd240 : gamma_data = 8'd253; 
	8'd241 : gamma_data = 8'd253; 
	8'd242 : gamma_data = 8'd253; 
	8'd243 : gamma_data = 8'd253; 
	8'd244 : gamma_data = 8'd254; 
	8'd245 : gamma_data = 8'd254; 
	8'd246 : gamma_data = 8'd254; 
	8'd247 : gamma_data = 8'd254; 
	8'd248 : gamma_data = 8'd254; 
	8'd249 : gamma_data = 8'd254; 
	8'd250 : gamma_data = 8'd254; 
	8'd251 : gamma_data = 8'd254; 
	8'd252 : gamma_data = 8'd255; 
	8'd253 : gamma_data = 8'd255; 
	8'd254 : gamma_data = 8'd255; 
	8'd255 : gamma_data = 8'd255; 
	endcase
end

endmodule
