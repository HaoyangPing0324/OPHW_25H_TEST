//�ӳ�1��ʱ���ź�
module binarization(

    input               clk             ,   
    input               rst_n           ,   
    input   [7:0]       y_in       ,

    output   [23:0]        data_bin            
);

//��һ���ÿ�����ֵ�����ַ�k��Ч�������䷱��������ÿ��ͼƬ��ֵ��һ��������Ǩ�ơ������Ҫ�ֲ���ֵ��
//parameter Binar_THRESHOLD = 128;
//parameter Binar_THRESHOLD = 192;
//parameter Binar_THRESHOLD = 160;
//parameter Binar_THRESHOLD = 144;
//parameter Binar_THRESHOLD = 152;
//parameter Binar_THRESHOLD = 156;
//parameter Binar_THRESHOLD = 158;
parameter Binar_THRESHOLD = 159;

reg pix;

//��ֵ��
always @(posedge clk or negedge rst_n) begin
    if(!rst_n)
        pix <= 1'b0;
    else if(y_in > Binar_THRESHOLD)  //��ֵ
        pix <= 1'b1;
    else
        pix <= 1'b0;
end

assign data_bin = {24{pix}};

endmodule 