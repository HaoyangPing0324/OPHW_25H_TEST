`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//Copyright(C) ����ԭ�� 2023-2033
// Revised By HaoyangPing_PKU
//
//////////////////////////////////////////////////////////////////////////////////
`define UD #1
module video_display # (
    parameter                            COCLOR_DEPP=8, // number of bits per channel
    parameter                            X_BITS=12,
    parameter                            Y_BITS=12,
    parameter                            H_ACT = 12'd1280,
    parameter                            V_ACT = 12'd720
)(                                       
    input                                rstn, 
    input                                pix_clk,
    input [X_BITS-1:0]                   act_x,
	input [Y_BITS-1:0]                   act_y,
    input                                vs_in, 
    input                                hs_in, 
    input                                de_in,
    
    output reg                           vs_out, 
    output reg                           hs_out, 
    output reg                           de_out,
    output reg [3*COCLOR_DEPP-1:0]       pixel_data 
);

    //parameter define     

localparam NUMBER_OF_DELAYED_CLKS = 3 ;//�ҶȻ��ӳ���3��ʱ���ź�
	
localparam PIC_WIDTH   = 12'd256;    //ͼƬ���
localparam PIC_HEIGHT  = 12'd256;    //ͼƬ�߶�
localparam PIC_X_START = 12'd640;     //ͼƬ��ʼ�������
localparam PIC_Y_START = 12'd412;     //ͼƬ��ʼ��������

localparam PIC_WIDTH2   = 12'd256;    //ͼƬ���
localparam PIC_HEIGHT2  = 12'd256;    //ͼƬ�߶�
localparam PIC_X_START2 = 12'd1024;     //ͼƬ��ʼ�������
localparam PIC_Y_START2 = 12'd412;     //ͼƬ��ʼ��������                       
                       
localparam BACK_COLOR  = 24'hE0FFFF; //����ɫ��ǳ��ɫ
//localparam BACK_COLOR  = 24'hFF0000; //����ɫ����ɫ�����Լ��������

//reg define
reg   [15:0]  rom_addr  ;  //ROM��ַ
reg   [15:0]  rom_addr1  ;  //ROM��ַ
reg   [15:0]  rom_addr2  ;  //ROM��ַ

//wire define   
wire  [23:0]  rom_rd_data ;//ROM����
wire  [23:0]  rom_rd_data2 ;//ROM����
wire vs_out0;
wire hs_out0;
wire de_out0;
wire [23:0] data_previous;
wire [23:0] data_after_process;

//*****************************************************
//**                    main code
//*****************************************************
//ΪLCD��ʾ�������ͼƬ
always @(posedge pix_clk or negedge rstn) begin
    if (!rstn)
        pixel_data <= BACK_COLOR;
    else if( (act_x >= PIC_X_START -1'b1) && (act_x < PIC_X_START + PIC_WIDTH -1'b1) 
          && (act_y >= PIC_Y_START) && (act_y < PIC_Y_START + PIC_HEIGHT) )
        pixel_data <= data_previous ;  //��ʾԭͼƬ
    else if( (act_x >= PIC_X_START2 -1'b1) && (act_x < PIC_X_START2 + PIC_WIDTH2 -1'b1) 
          && (act_y >= PIC_Y_START2) && (act_y < PIC_Y_START2 + PIC_HEIGHT2) )
        pixel_data <= data_after_process ;  //��ʾ�����ͼƬ
    else
        pixel_data <= BACK_COLOR;        //��Ļ����ɫ
end

always @(posedge pix_clk or negedge rstn) begin
    if (!rstn)
        rom_addr <= 16'd0;
    else if( (act_x >= PIC_X_START -2'd2 - NUMBER_OF_DELAYED_CLKS ) && (act_x < PIC_X_START + PIC_WIDTH -2'd2 - NUMBER_OF_DELAYED_CLKS ) 
          && (act_y >= PIC_Y_START) && (act_y < PIC_Y_START + PIC_HEIGHT) )
        rom_addr <= rom_addr1;  //��ʾԭͼƬ
    else if( (act_x >= PIC_X_START2 -2'd2 - NUMBER_OF_DELAYED_CLKS ) && (act_x < PIC_X_START2 + PIC_WIDTH2 -2'd2 - NUMBER_OF_DELAYED_CLKS ) 
          && (act_y >= PIC_Y_START2) && (act_y < PIC_Y_START2 + PIC_HEIGHT2) )
        rom_addr <= rom_addr2;  //��ʾ�����ͼƬ
    else
        rom_addr <= 16'd0;        //��Ļ����ɫ
end

//���ݵ�ǰɨ���ĺ�������ΪROM��ַ��ֵ
always @(posedge pix_clk or negedge rstn) begin
    if(!rstn)
        rom_addr1 <= 16'd0;
    //����������λ��ͼƬ��ʾ����ʱ,�ۼ�ROM��ַ    
    else if( (act_x >= PIC_X_START -2'd2 - NUMBER_OF_DELAYED_CLKS ) && (act_x < PIC_X_START + PIC_WIDTH -2'd2 - NUMBER_OF_DELAYED_CLKS ) 
          && (act_y >= PIC_Y_START) && (act_y < PIC_Y_START + PIC_HEIGHT) )
        rom_addr1 <= rom_addr1 + 1'b1;
    //����������λ��ͼƬ�������һ�����ص�ʱ,ROM��ַ����    
    else if((act_y >= PIC_Y_START + PIC_HEIGHT))
        rom_addr1 <= 16'd0;
end

always @(posedge pix_clk or negedge rstn) begin
    if(!rstn)
        rom_addr2 <= 16'd0;
    //����������λ��ͼƬ��ʾ����ʱ,�ۼ�ROM��ַ    
    else if( (act_x >= PIC_X_START2 -2'd2 - NUMBER_OF_DELAYED_CLKS ) && (act_x < PIC_X_START2 + PIC_WIDTH2 -2'd2 - NUMBER_OF_DELAYED_CLKS ) 
          && (act_y >= PIC_Y_START2) && (act_y < PIC_Y_START2 + PIC_HEIGHT2) )
        rom_addr2 <= rom_addr2 + 1'b1;
    //����������λ��ͼƬ�������һ�����ص�ʱ,ROM��ַ����    
    else if((act_y >= PIC_Y_START + PIC_HEIGHT))
        rom_addr2 <= 16'd0;
end



//ROM���洢ͼƬ
blk_mem_gen_0 blk_mem_gen_0 (
  .addr    (rom_addr),          // input [15:0]
  .clk     (pix_clk),          // input
  .rst     (~rstn),            // input
  .rd_data (rom_rd_data)     	// output [23:0]
);

//ͼƬ����
RGB2YCbCr u_RGB2YCbCr (
    .clk          (pix_clk),           // ���룺ģ��ʱ��
    .rst_n        (rstn),         // ���룺�첽��λ���͵�ƽ��Ч
    .img_data_in  (rom_rd_data),   // ���룺24λRGB�������� [23:0]
    .data_ycbcr   (data_after_process) // �����24λYCbCr������� [23:0]
);


// ʵ����ͬ���ź��ӳ�ģ��
signal_delay #(
    .NUMBER_OF_DELAYED_CLKS (NUMBER_OF_DELAYED_CLKS)
) u_signal_delay (
    .rstn     (rstn),
    .clk      (pix_clk),
    .vs_in    (vs_in),
    .hs_in    (hs_in),
    .de_in    (de_in),
    .vs_out   (vs_out0),
    .hs_out   (hs_out0),
    .de_out   (de_out0)
);

    always @(posedge pix_clk)//��ģ���Դ���һ��ʱ���ӳ�
    begin
        vs_out <= `UD vs_out0;
        hs_out <= `UD hs_out0;
        de_out <= `UD de_out0;
    end

// ʵ���������ź��ӳ�ģ��
data_delay #(
    .NUMBER_OF_DELAYED_CLKS (NUMBER_OF_DELAYED_CLKS),
    .COCLOR_DEPP            (COCLOR_DEPP)
) u_data_delay (
    .rstn     (rstn),
    .clk      (pix_clk),
    .data_in  (rom_rd_data),
    .data_out (data_previous)
);

endmodule
