`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//Author: HaoyangPing_PKU
//////////////////////////////////////////////////////////////////////////////////
`define UD #1
module video_display # (
    parameter                            COCLOR_DEPP=8, // number of bits per channel
    parameter                            X_BITS=12,
    parameter                            Y_BITS=12,
    parameter                            H_ACT = 12'd1280,
    parameter                            V_ACT = 12'd720
)(                                       
    input                                rstn, 
    input                                pix_clk,
    input [X_BITS-1:0]                   act_x,
	input [Y_BITS-1:0]                   act_y,
    input                                vs_in, 
    input                                hs_in, 
    input                                de_in,
    
    output reg                           vs_out, 
    output reg                           hs_out, 
    output reg                           de_out,
    output reg [3*COCLOR_DEPP-1:0]       pixel_data 
);

//parameter define     
//��˹�˲� 4+2clks
localparam NUMBER_OF_DELAYED_CLKS_PREVIOUS = 6 ;

localparam PIC_WIDTH   = 12'd256;    //ͼƬ���
localparam PIC_HEIGHT  = 12'd256;    //ͼƬ�߶�

localparam PIC_X_START_COL1 = 12'd640;     //ͼƬ��ʼ�������
localparam PIC_X_START_COL2 = 12'd1024;

localparam PIC_Y_START_ROW = 12'd412;     //ͼƬ��ʼ��������                   
                       
localparam BACK_COLOR  = 24'hE0FFFF; //����ɫ��ǳ��ɫ
//localparam BACK_COLOR  = 24'hFF0000; //����ɫ����ɫ�����Լ��������

//reg define
reg   [15:0]  rom_addr  ;  //ROM��ַ
reg [15:0] rom_addr_previous;
reg [15:0] rom_addr_gauss_filter;

//wire define
wire vs_out0;
wire hs_out0;
wire de_out0;  

wire  [23:0]  rom_rd_data ;//ROM����

wire [23:0] data_previous;

wire [23:0] data_gauss_filter;

wire [7:0] matrix11[0:2];
wire [7:0] matrix12[0:2];
wire [7:0] matrix13[0:2];
wire [7:0] matrix21[0:2];
wire [7:0] matrix22[0:2];
wire [7:0] matrix23[0:2];
wire [7:0] matrix31[0:2];
wire [7:0] matrix32[0:2];
wire [7:0] matrix33[0:2];

//*****************************************************
//**                    main code
//*****************************************************
//ΪLCD��ʾ�������ͼƬ
always @(posedge pix_clk or negedge rstn) begin
    if (!rstn)
        pixel_data <= BACK_COLOR;
    else if( (act_x >= PIC_X_START_COL1 -1'b1) && (act_x < PIC_X_START_COL1 + PIC_WIDTH -1'b1) 
          && (act_y >= PIC_Y_START_ROW) && (act_y < PIC_Y_START_ROW + PIC_HEIGHT) )
        pixel_data <= data_previous ;  //��ʾԭͼƬ
	else if( (act_x >= PIC_X_START_COL2 -1'b1) && (act_x < PIC_X_START_COL2 + PIC_WIDTH -1'b1) 
          && (act_y >= PIC_Y_START_ROW) && (act_y < PIC_Y_START_ROW + PIC_HEIGHT) )
        pixel_data <= data_gauss_filter ;  //��ʾ��˹�˲�ͼƬ
    else
        pixel_data <= BACK_COLOR;        //��Ļ����ɫ
end


always @(posedge pix_clk or negedge rstn) begin
    if (!rstn)
        rom_addr <= 16'd0;		
	else if( (act_x >= PIC_X_START_COL1 -2'd2 -NUMBER_OF_DELAYED_CLKS_PREVIOUS) && (act_x < PIC_X_START_COL1 + PIC_WIDTH -2'd2 -NUMBER_OF_DELAYED_CLKS_PREVIOUS) 
		&& (act_y >= PIC_Y_START_ROW) && (act_y < PIC_Y_START_ROW + PIC_HEIGHT) )//��ʾԭͼƬ
        rom_addr <= rom_addr_previous;
    else if( (act_x >= PIC_X_START_COL2 -2'd2 -NUMBER_OF_DELAYED_CLKS_PREVIOUS) && (act_x < PIC_X_START_COL2 + PIC_WIDTH -2'd2 -NUMBER_OF_DELAYED_CLKS_PREVIOUS) 
		&& (act_y >= PIC_Y_START_ROW) && (act_y < PIC_Y_START_ROW + PIC_HEIGHT) )//��ʾ��˹�˲�ͼƬ
        rom_addr <= rom_addr_gauss_filter; 
    else
        rom_addr <= 16'd0;        //��Ļ����ɫ
end

//���ݵ�ǰɨ���ĺ�������ΪROM��ַ��ֵ
always @(posedge pix_clk or negedge rstn) begin
    if(!rstn)
        rom_addr_previous <= 16'd0;
    // ����������λ��ͼƬ��ʾ����ʱ,�ۼ�ROM��ַ
    else if( (act_x >= PIC_X_START_COL1 - 2'd2 - NUMBER_OF_DELAYED_CLKS_PREVIOUS) && 
             (act_x < PIC_X_START_COL1 + PIC_WIDTH - 2'd2 - NUMBER_OF_DELAYED_CLKS_PREVIOUS) && 
             (act_y >= PIC_Y_START_ROW) && 
             (act_y < PIC_Y_START_ROW + PIC_HEIGHT) )
        rom_addr_previous <= rom_addr_previous + 1'b1;
    // ����������λ��ͼƬ�������һ�����ص�ʱ,ROM��ַ����
    else if((act_y >= PIC_Y_START_ROW + PIC_HEIGHT))
        rom_addr_previous <= 16'd0;
end

always @(posedge pix_clk or negedge rstn) begin
    if(!rstn)
        rom_addr_gauss_filter <= 16'd0;
    // ����������λ��ͼƬ��ʾ����ʱ,�ۼ�ROM��ַ
    else if( (act_x >= PIC_X_START_COL2 - 2'd2 - NUMBER_OF_DELAYED_CLKS_PREVIOUS) && 
             (act_x < PIC_X_START_COL2 + PIC_WIDTH - 2'd2 - NUMBER_OF_DELAYED_CLKS_PREVIOUS) && 
             (act_y >= PIC_Y_START_ROW) && 
             (act_y < PIC_Y_START_ROW + PIC_HEIGHT) )
        rom_addr_gauss_filter <= rom_addr_gauss_filter + 1'b1;
    // ����������λ��ͼƬ�������һ�����ص�ʱ,ROM��ַ����
    else if((act_y >= PIC_Y_START_ROW + PIC_HEIGHT))
        rom_addr_gauss_filter <= 16'd0;
end

//ROM���洢ͼƬ
blk_mem_gen_0 blk_mem_gen_0 (
  .addr    (rom_addr),          // input [15:0]
  .clk     (pix_clk),          // input
  .rst     (~rstn),            // input
  .rd_data (rom_rd_data)     	// output [23:0]
);

//ͼƬ����
//��˹�˲�

genvar i;
generate
    for (i = 0; i <= 2; i = i + 1) begin : u_data_gauss_filter
        matrix_3x3 
		#(
			.IMG_WIDTH (12'd2200),
			.IMG_HEIGHT(12'd1125)
		)
		u_matrix_3x3
		(
			.video_clk  (pix_clk),
			.rst_n      (rstn),
			.video_data (rom_rd_data[(23 - 8 *i):(16 - 8*i)]),
			.matrix11   (matrix11[i]),
			.matrix12   (matrix12[i]),
			.matrix13   (matrix13[i]),
			.matrix21   (matrix21[i]),
			.matrix22   (matrix22[i]),
			.matrix23   (matrix23[i]),
			.matrix31   (matrix31[i]),
			.matrix32   (matrix32[i]),
			.matrix33   (matrix33[i])
		);
		
		gauss_filter u_gauss_filter
		(
			.video_clk        (pix_clk),        // ������Ƶʱ��
			.rst_n            (rstn),            // ��λ�źţ��͵�ƽ��Ч
    
			// 3x3������������
			.matrix11         (matrix11[i]),         // ��1�е�1������
			.matrix12         (matrix12[i]),         // ��1�е�2������  
			.matrix13         (matrix13[i]),         // ��1�е�3������
			.matrix21         (matrix21[i]),         // ��2�е�1������
			.matrix22         (matrix22[i]),         // ��2�е�2������
			.matrix23         (matrix23[i]),         // ��2�е�3������
			.matrix31         (matrix31[i]),         // ��3�е�1������
			.matrix32         (matrix32[i]),         // ��3�е�2������
			.matrix33         (matrix33[i]),         // ��3�е�3������
		
			.gauss_filter_data (data_gauss_filter[(23 - 8 *i):(16 - 8*i)])  // ��˹�˲��������
		);
    end
endgenerate

// ʵ����ͬ���ź��ӳ�ģ��
signal_delay #(
    .NUMBER_OF_DELAYED_CLKS (NUMBER_OF_DELAYED_CLKS_PREVIOUS)
) u_signal_delay (
    .rstn     (rstn),
    .clk      (pix_clk),
    .vs_in    (vs_in),
    .hs_in    (hs_in),
    .de_in    (de_in),
    .vs_out   (vs_out0),
    .hs_out   (hs_out0),
    .de_out   (de_out0)
);

    always @(posedge pix_clk)//��ģ���Դ���һ��ʱ���ӳ�
    begin
        vs_out <= `UD vs_out0;
        hs_out <= `UD hs_out0;
        de_out <= `UD de_out0;
    end

// ʵ���������ź��ӳ�ģ��
data_delay #(
            .NUMBER_OF_DELAYED_CLKS (NUMBER_OF_DELAYED_CLKS_PREVIOUS),
            .COCLOR_DEPP            (COCLOR_DEPP)
        ) u_data_delay_inst (
            .rstn     (rstn),
            .clk      (pix_clk),
            .data_in  (rom_rd_data),
            .data_out (data_previous)
);

endmodule
