module rom_test_top
(
    input    wire               rd_clk        ,//��ʱ��
    input    wire               rst_n         ,//��λ



    input    wire    [9:0]      rd_addr       ,//����ַ

    
    output   wire    [63:0]      rd_data        //������
    
   
);


rom_test rom_test_inst (
  .addr(rd_addr),          // input [9:0]
  .clk(rd_clk),            // input
  .rst(~rst_n),            // input
  .rd_data(rd_data)     // output [63:0]
);




endmodule