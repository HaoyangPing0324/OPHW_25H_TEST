module ram_test_top
(
    input    wire               wr_clk        ,//дʱ��
    input    wire               rd_clk        ,//��ʱ��
    input    wire               rst_n         ,//��λ

    input    wire               rw_en         ,//��дʹ���ź�
    input    wire    [5:0]      wr_addr       ,//д��ַ
    input    wire    [5:0]      rd_addr       ,//����ַ
    input    wire    [7:0]      wr_data       ,//д����
    
    output   wire    [7:0]      rd_data        //������
);


ram_test ram_test_inst (
  .wr_data(wr_data),    // input [7:0]
  .wr_addr(wr_addr),    // input [5:0]
  .wr_en(rw_en),        // input    
  .wr_clk(wr_clk),      // input
  .wr_rst(~rst_n),      // input

  .rd_addr(rd_addr),    // input [5:0]
  .rd_data(rd_data),    // output [7:0]
  .rd_clk(rd_clk),      // input
  .rd_rst(~rst_n)       // input
);



endmodule