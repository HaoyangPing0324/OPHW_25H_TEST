`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//Author: HaoyangPing_PKU
//////////////////////////////////////////////////////////////////////////////////
`define UD #1
module video_display # (
    parameter                            COCLOR_DEPP=8, // number of bits per channel
    parameter                            X_BITS=12,
    parameter                            Y_BITS=12,
    parameter                            H_ACT = 12'd1280,
    parameter                            V_ACT = 12'd720
)(                                       
    input                                rstn, 
    input                                pix_clk,
    input [X_BITS-1:0]                   act_x,
	input [Y_BITS-1:0]                   act_y,
    input                                vs_in, 
    input                                hs_in, 
    input                                de_in,
    
    output reg                           vs_out, 
    output reg                           hs_out, 
    output reg                           de_out,
    output reg [3*COCLOR_DEPP-1:0]       pixel_data 
);

    //parameter define     
//�ҶȻ� 3 clk
//��ֵ�� 3+1 clk
//�ֲ���ֵ�� 3+6 clk
localparam NUMBER_OF_DELAYED_CLKS_PREVIOUS = 9 ;
localparam NUMBER_OF_DELAYED_CLKS_GREY = 6 ;
localparam NUMBER_OF_DELAYED_CLKS_BIN = 5 ;
	
localparam PIC_WIDTH   = 12'd256;    //ͼƬ���
localparam PIC_HEIGHT  = 12'd256;    //ͼƬ�߶�
localparam PIC_X_START = 12'd256;     //ͼƬ��ʼ�������
localparam PIC_Y_START = 12'd412;     //ͼƬ��ʼ��������

localparam PIC_WIDTH_GREY   = 12'd256;    //ͼƬ���
localparam PIC_HEIGHT_GREY  = 12'd256;    //ͼƬ�߶�
localparam PIC_X_START_GREY = 12'd640;     //ͼƬ��ʼ�������
localparam PIC_Y_START_GREY = 12'd412;     //ͼƬ��ʼ��������

localparam PIC_WIDTH_BIN   = 12'd256;    //ͼƬ���
localparam PIC_HEIGHT_BIN  = 12'd256;    //ͼƬ�߶�
localparam PIC_X_START_BIN = 12'd1024;     //ͼƬ��ʼ�������
localparam PIC_Y_START_BIN = 12'd412;     //ͼƬ��ʼ�������� 

localparam PIC_WIDTH_AREA_BIN   = 12'd256;    //ͼƬ���
localparam PIC_HEIGHT_AREA_BIN  = 12'd256;    //ͼƬ�߶�
//localparam PIC_X_START_AREA_BIN = 12'd10;     //ͼƬ��ʼ�������
//localparam PIC_Y_START_AREA_BIN = 12'd10;     //ͼƬ��ʼ�������� 
localparam PIC_X_START_AREA_BIN = 12'd1408;     //ͼƬ��ʼ�������
localparam PIC_Y_START_AREA_BIN = 12'd412;     //ͼƬ��ʼ�������� 
                       
                       
localparam BACK_COLOR  = 24'hE0FFFF; //����ɫ��ǳ��ɫ
//localparam BACK_COLOR  = 24'hFF0000; //����ɫ����ɫ�����Լ��������

//reg define
reg   [15:0]  rom_addr  ;  //ROM��ַ
reg   [15:0]  rom_addr_previous  ;  //ROM��ַ
reg   [15:0]  rom_addr_grey  ;  //ROM��ַ
reg   [15:0]  rom_addr_bin  ;  //ROM��ַ
reg   [15:0]  rom_addr_area_bin  ;  //ROM��ַ

//wire define 
wire vs_out0;
wire hs_out0;
wire de_out0;  

wire  [23:0]  rom_rd_data ;//ROM����

wire [23:0] data_previous;
wire [23:0] data_after_grey;
wire [23:0] data_after_bin;
wire [23:0] data_after_grey_d;
wire [23:0] data_after_bin_d;
wire [23:0] data_after_area_bin;



//*****************************************************
//**                    main code
//*****************************************************
//ΪLCD��ʾ�������ͼƬ
always @(posedge pix_clk or negedge rstn) begin
    if (!rstn)
        pixel_data <= BACK_COLOR;
    else if( (act_x >= PIC_X_START -1'b1) && (act_x < PIC_X_START + PIC_WIDTH -1'b1) 
          && (act_y >= PIC_Y_START) && (act_y < PIC_Y_START + PIC_HEIGHT) )
        pixel_data <= data_previous ;  //��ʾԭͼƬ
    else if( (act_x >= PIC_X_START_GREY -1'b1) && (act_x < PIC_X_START_GREY + PIC_WIDTH_GREY -1'b1) 
          && (act_y >= PIC_Y_START_GREY) && (act_y < PIC_Y_START_GREY + PIC_HEIGHT_GREY) )
        pixel_data <= data_after_grey_d ;  //�ҶȻ���ͼƬ
    else if( (act_x >= PIC_X_START_BIN -1'b1) && (act_x < PIC_X_START_BIN + PIC_WIDTH_BIN -1'b1) 
          && (act_y >= PIC_Y_START_BIN) && (act_y < PIC_Y_START_BIN + PIC_HEIGHT_BIN) )
        pixel_data <= data_after_bin_d ;  //��ֵ����ͼƬ
    else if( (act_x >= PIC_X_START_AREA_BIN -1'b1) && (act_x < PIC_X_START_AREA_BIN + PIC_WIDTH_AREA_BIN -1'b1) 
          && (act_y >= PIC_Y_START_AREA_BIN) && (act_y < PIC_Y_START_AREA_BIN + PIC_HEIGHT_AREA_BIN) )
        //pixel_data <= data_after_bin_d ;  //��ֵ����ͼƬ
        pixel_data <= data_after_area_bin ;  //�ֲ���ֵ����ͼƬ
    else
        pixel_data <= BACK_COLOR;        //��Ļ����ɫ
//������
//pixel_data <= data_after_area_bin ;  //�ֲ���ֵ����ͼƬ
end

always @(posedge pix_clk or negedge rstn) begin
    if (!rstn)
        rom_addr <= 16'd0;
    else if( (act_x >= PIC_X_START -2'd2 -NUMBER_OF_DELAYED_CLKS_PREVIOUS ) && (act_x < PIC_X_START + PIC_WIDTH -2'd2 -NUMBER_OF_DELAYED_CLKS_PREVIOUS) 
          && (act_y >= PIC_Y_START) && (act_y < PIC_Y_START + PIC_HEIGHT) )
        rom_addr <= rom_addr_previous;  //��ʾԭͼƬ
    else if( (act_x >= PIC_X_START_GREY -2'd2 - NUMBER_OF_DELAYED_CLKS_PREVIOUS) && (act_x < PIC_X_START_GREY + PIC_WIDTH_GREY  -2'd2 -NUMBER_OF_DELAYED_CLKS_PREVIOUS) 
          && (act_y >= PIC_Y_START_GREY) && (act_y < PIC_Y_START_GREY + PIC_HEIGHT_GREY) )
        rom_addr <= rom_addr_grey;  //�ҶȻ���ͼƬ
    else if( (act_x >= PIC_X_START_BIN -2'd2 - NUMBER_OF_DELAYED_CLKS_PREVIOUS ) && (act_x < PIC_X_START_BIN + PIC_WIDTH_BIN -2'd2 -NUMBER_OF_DELAYED_CLKS_PREVIOUS) 
          && (act_y >= PIC_Y_START_BIN) && (act_y < PIC_Y_START_BIN + PIC_HEIGHT_BIN) )
        rom_addr <= rom_addr_bin;  //��ֵ����ͼƬ
    else if( (act_x >= PIC_X_START_AREA_BIN -2'd2 -NUMBER_OF_DELAYED_CLKS_PREVIOUS) && (act_x < PIC_X_START_AREA_BIN + PIC_WIDTH_AREA_BIN --2'd2 -NUMBER_OF_DELAYED_CLKS_PREVIOUS) 
          && (act_y >= PIC_Y_START_AREA_BIN) && (act_y < PIC_Y_START_AREA_BIN + PIC_HEIGHT_AREA_BIN) )
        rom_addr <= rom_addr_area_bin;  //�ֲ���ֵ����ͼƬ
    else
        rom_addr <= 16'd0;        //��Ļ����ɫ
end

//���ݵ�ǰɨ���ĺ�������ΪROM��ַ��ֵ
always @(posedge pix_clk or negedge rstn) begin
    if(!rstn)
        rom_addr_previous <= 16'd0;
    //����������λ��ͼƬ��ʾ����ʱ,�ۼ�ROM��ַ    
    else if( (act_x >= PIC_X_START -2'd2 -NUMBER_OF_DELAYED_CLKS_PREVIOUS ) && (act_x < PIC_X_START + PIC_WIDTH -2'd2 -NUMBER_OF_DELAYED_CLKS_PREVIOUS) 
          && (act_y >= PIC_Y_START) && (act_y < PIC_Y_START + PIC_HEIGHT) )
        rom_addr_previous <= rom_addr_previous + 1'b1;
    //����������λ��ͼƬ�������һ�����ص�ʱ,ROM��ַ����    
    else if((act_y >= PIC_Y_START + PIC_HEIGHT))
        rom_addr_previous <= 16'd0;
end

always @(posedge pix_clk or negedge rstn) begin
    if(!rstn)
        rom_addr_grey <= 16'd0;
    //����������λ��ͼƬ��ʾ����ʱ,�ۼ�ROM��ַ    
   else if( (act_x >= PIC_X_START_GREY -2'd2 -NUMBER_OF_DELAYED_CLKS_PREVIOUS) && (act_x < PIC_X_START_GREY + PIC_WIDTH_GREY -2'd2 -NUMBER_OF_DELAYED_CLKS_PREVIOUS) 
          && (act_y >= PIC_Y_START_GREY) && (act_y < PIC_Y_START_GREY + PIC_HEIGHT_GREY) )
        rom_addr_grey <= rom_addr_grey + 1'b1;
    //����������λ��ͼƬ�������һ�����ص�ʱ,ROM��ַ����    
    else if((act_y >= PIC_Y_START + PIC_HEIGHT))
        rom_addr_grey <= 16'd0;
end

always @(posedge pix_clk or negedge rstn) begin
    if(!rstn)
        rom_addr_bin <= 16'd0;
    //����������λ��ͼƬ��ʾ����ʱ,�ۼ�ROM��ַ    
   else if( (act_x >= PIC_X_START_BIN -2'd2 -NUMBER_OF_DELAYED_CLKS_PREVIOUS) && (act_x < PIC_X_START_BIN + PIC_WIDTH_BIN -2'd2 -NUMBER_OF_DELAYED_CLKS_PREVIOUS) 
          && (act_y >= PIC_Y_START_BIN) && (act_y < PIC_Y_START_BIN + PIC_HEIGHT_BIN) )
        rom_addr_bin <= rom_addr_bin + 1'b1;
    //����������λ��ͼƬ�������һ�����ص�ʱ,ROM��ַ����    
    else if((act_y >= PIC_Y_START + PIC_HEIGHT))
        rom_addr_bin <= 16'd0;
end

always @(posedge pix_clk or negedge rstn) begin
    if(!rstn)
        rom_addr_area_bin <= 16'd0;
    //����������λ��ͼƬ��ʾ����ʱ,�ۼ�ROM��ַ    
   else if( (act_x >= PIC_X_START_AREA_BIN -2'd2 -NUMBER_OF_DELAYED_CLKS_PREVIOUS) && (act_x < PIC_X_START_AREA_BIN + PIC_WIDTH_AREA_BIN -2'd2 -NUMBER_OF_DELAYED_CLKS_PREVIOUS) 
          && (act_y >= PIC_Y_START_AREA_BIN) && (act_y < PIC_Y_START_AREA_BIN + PIC_HEIGHT_AREA_BIN) )
        rom_addr_area_bin <= rom_addr_area_bin + 1'b1;
    //����������λ��ͼƬ�������һ�����ص�ʱ,ROM��ַ����    
    else if((act_y >= PIC_Y_START + PIC_HEIGHT))
        rom_addr_area_bin <= 16'd0;
end

//ROM���洢ͼƬ
blk_mem_gen_0 blk_mem_gen_0 (
  .addr    (rom_addr),          // input [15:0]
  .clk     (pix_clk),          // input
  .rst     (~rstn),            // input
  .rd_data (rom_rd_data)     	// output [23:0]
);

//ͼƬ����
//�ҶȻ�
RGB2YCbCr u_RGB2YCbCr (
    .clk          (pix_clk),           // ���룺ģ��ʱ��
    .rst_n        (rstn),         // ���룺�첽��λ���͵�ƽ��Ч
    .img_data_in  (rom_rd_data),   // ���룺24λRGB�������� [23:0]
    .data_ycbcr   (data_after_grey) // �����24λYCbCr������� [23:0]
);

//��ֵ��
binarization u_binarization (
    .clk     (pix_clk),          // ���룺ʱ���ź�
    .rst_n   (rstn),        // ���룺�첽��λ���͵�ƽ��Ч
    .y_in    (data_after_grey[7:0]),    // ���룺8λY�������� [7:0]
    .data_bin     (data_after_bin)    // �������ֵ�����ؽ��
);

//�ֲ���ֵ��
area_bin#(
    	.IMG_WIDTH(12'd2200)	,
		.IMG_HEIGHT(12'd1125)
)u_area_bin
(
    .video_clk      (pix_clk),     // ���룺��Ƶʱ��
    .rst_n          (rstn),         // ���룺�첽��λ���͵�ƽ��Ч
    .video_data (data_after_grey[7:0]),  // ���룺8λ�������� [7:0]
    
    .data_area_bin  (data_after_area_bin) // ����������ֵ�����
);

// ʵ����ͬ���ź��ӳ�ģ��
signal_delay #(
    .NUMBER_OF_DELAYED_CLKS (NUMBER_OF_DELAYED_CLKS_PREVIOUS)
) u_signal_delay (
    .rstn     (rstn),
    .clk      (pix_clk),
    .vs_in    (vs_in),
    .hs_in    (hs_in),
    .de_in    (de_in),
    .vs_out   (vs_out0),
    .hs_out   (hs_out0),
    .de_out   (de_out0)
);

    always @(posedge pix_clk)//��ģ���Դ���һ��ʱ���ӳ�
    begin
        vs_out <= `UD vs_out0;
        hs_out <= `UD hs_out0;
        de_out <= `UD de_out0;
    end

// ʵ���������ź��ӳ�ģ��
data_delay #(
    .NUMBER_OF_DELAYED_CLKS (NUMBER_OF_DELAYED_CLKS_PREVIOUS),
    .COCLOR_DEPP            (COCLOR_DEPP)
) u_data_delay_previous (
    .rstn     (rstn),
    .clk      (pix_clk),
    .data_in  (rom_rd_data),
    .data_out (data_previous)
);

data_delay #(
    .NUMBER_OF_DELAYED_CLKS (NUMBER_OF_DELAYED_CLKS_GREY),
    .COCLOR_DEPP            (COCLOR_DEPP)
) u_data_delay_grey (
    .rstn     (rstn),
    .clk      (pix_clk),
    .data_in  (data_after_grey),
    .data_out (data_after_grey_d)
);

data_delay #(
    .NUMBER_OF_DELAYED_CLKS (NUMBER_OF_DELAYED_CLKS_BIN),
    .COCLOR_DEPP            (COCLOR_DEPP)
) u_data_delay_bin (
    .rstn     (rstn),
    .clk      (pix_clk),
    .data_in  (data_after_bin),
    .data_out (data_after_bin_d)
);
endmodule
